module hazard_det_unit (
    
);

endmodule