module immediate_gen (
    input  wire [31:0] instr,
    output reg  [63:0] imm_out
);
    
endmodule
