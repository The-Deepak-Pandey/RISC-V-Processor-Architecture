`include "control.v"
`include "register_file.v"
`include "immediate_gen.v"

module instruction_decode_stage(
    intput wire 
);

endmodule