module seq_processor(
    input wire clk,
    input wire rst;
);

    

endmodule