module write_back(
    input mem_read,
    input [4:0] rd_addr,
    input [63:0] mem_data,
    output reg [63:0] write_data,
);

    

endmodule